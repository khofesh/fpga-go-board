module VGA_Test_Patterns_Top (
    input i_Clk, // main clock
    input i_UART_RX, // uart rx data
    output o_UART_TX, // uart tx data
    // segment1 is upper digit, segment2 is lower digit
    output o_Segment1_A,
    output o_Segment1_B,
    output o_Segment1_C,
    output o_Segment1_D,
    output o_Segment1_E,
    output o_Segment1_F,
    output o_Segment1_G,
    // 
    output o_Segment2_A,
    output o_Segment2_B,
    output o_Segment2_C,
    output o_Segment2_D,
    output o_Segment2_E,
    output o_Segment2_F,
    output o_Segment2_G,

    // vga
    output o_VGA_HSync,
    output o_VGA_VSync,
    output o_VGA_Red_0,
    output o_VGA_Red_1,
    output o_VGA_Grn_0,
    output o_VGA_Grn_1,
    output o_VGA_Grn_2,
    output o_VGA_Blu_0,
    output o_VGA_Blu_1,
    output o_VGA_Blu_2
);

    // vga constants to set frame size
    parameter c_VIDEO_WIDTH = 3;
    parameter c_TOTAL_COLS = 800;
    parameter c_TOTAL_ROWS = 525;
    parameter c_ACTIVE_COLS = 640;
    parameter c_ACTIVE_ROWS = 480;

    wire w_RX_DV;
    wire [7:0] w_RX_Byte;
    wire w_TX_Active, w_TX_Serial;
    
    wire w_Segment1_A, w_Segment2_A;
    wire w_Segment1_B, w_Segment2_B;
    wire w_Segment1_C, w_Segment2_C;
    wire w_Segment1_D, w_Segment2_D;
    wire w_Segment1_E, w_Segment2_E;
    wire w_Segment1_F, w_Segment2_F;
    wire w_Segment1_G, w_Segment2_G;

    reg [3:0] r_TP_Index = 0;

    // common vga signals
    wire [c_VIDEO_WIDTH-1:0] w_Red_Video_TP, w_Red_Video_Porch;
    wire [c_VIDEO_WIDTH-1:0] w_Grn_Video_TP, w_Grn_Video_Porch;
    wire [c_VIDEO_WIDTH-1:0] w_Blu_Video_TP, w_Blu_Video_Porch;

    // 25,000,000 / 115,200 = 217
    UART_RX #(.CLKS_PER_BIT(217)) UART_RX_Inst
    (.i_Clock(i_Clk),
    .i_RX_Serial(i_UART_RX),
    .o_RX_DV(w_RX_DV),
    .o_RX_Byte(w_RX_Byte));

    UART_TX #(.CLKS_PER_BIT(217)) UART_TX_Inst
    (.i_Clock(i_Clk),
    .i_TX_DV(w_RX_DV), // pass rx to tx module for loopback
    .i_TX_Byte(w_RX_Byte), // pass rx to tx module for loopback
    .o_TX_Active(w_TX_Active),
    .o_TX_Serial(w_TX_Serial),
    .o_TX_Done());

    // drive UART line high when transmitter is not active
    assign o_UART_TX = w_TX_Active ? w_TX_Serial : 1'b1;

    // binary to 7-segment converter for upper digit
    Binary_To_7Segment SevenSeg1_Inst
    (.i_Clk(i_Clk),
     .i_Binary_Num(w_RX_Byte[7:4]),
     .o_Segment_A(w_Segment1_A),
     .o_Segment_B(w_Segment1_B),
     .o_Segment_C(w_Segment1_C),
     .o_Segment_D(w_Segment1_D),
     .o_Segment_E(w_Segment1_E),
     .o_Segment_F(w_Segment1_F),
     .o_Segment_G(w_Segment1_G));
    
    assign o_Segment1_A = ~w_Segment1_A;
    assign o_Segment1_B = ~w_Segment1_B;
    assign o_Segment1_C = ~w_Segment1_C;
    assign o_Segment1_D = ~w_Segment1_D;
    assign o_Segment1_E = ~w_Segment1_E;
    assign o_Segment1_F = ~w_Segment1_F;
    assign o_Segment1_G = ~w_Segment1_G;
    
    
    // Binary to 7-Segment Converter for Lower Digit
    Binary_To_7Segment SevenSeg2_Inst
    (.i_Clk(i_Clk),
     .i_Binary_Num(w_RX_Byte[3:0]),
     .o_Segment_A(w_Segment2_A),
     .o_Segment_B(w_Segment2_B),
     .o_Segment_C(w_Segment2_C),
     .o_Segment_D(w_Segment2_D),
     .o_Segment_E(w_Segment2_E),
     .o_Segment_F(w_Segment2_F),
     .o_Segment_G(w_Segment2_G));
    
    assign o_Segment2_A = ~w_Segment2_A;
    assign o_Segment2_B = ~w_Segment2_B;
    assign o_Segment2_C = ~w_Segment2_C;
    assign o_Segment2_D = ~w_Segment2_D;
    assign o_Segment2_E = ~w_Segment2_E;
    assign o_Segment2_F = ~w_Segment2_F;
    assign o_Segment2_G = ~w_Segment2_G;

    always @(posedge i_Clk) begin
        if (w_RX_DV == 1'b1) begin
            r_TP_Index <= w_RX_Byte[3:0];
        end
    end

    // generates sync pulses to run VGA
    VGA_Sync_Pulses #(.TOTAL_COLS(c_TOTAL_COLS),
        .TOTAL_ROWS(c_TOTAL_ROWS),
        .ACTIVE_COLS(c_ACTIVE_COLS),
        .ACTIVE_ROWS(c_ACTIVE_ROWS)) VGA_Sync_Pulses_Inst
    (.i_Clk(i_Clk),
    .o_HSync(w_HSync_Start),
    .o_VSync(w_VSync_Start),
    .o_Col_Count(),
    .o_Row_Count()
    );

    // drives red/green/blue video - test pattern 5 (color bars)
    Test_Pattern_Gen #(.VIDEO_WIDTH(c_VIDEO_WIDTH),
        .TOTAL_COLS(c_TOTAL_COLS),
        .TOTAL_ROWS(c_TOTAL_ROWS),
        .ACTIVE_COLS(c_ACTIVE_COLS),
        .ACTIVE_ROWS(c_ACTIVE_ROWS))
    Test_Pattern_Gen_Inst
    (.i_Clk(i_Clk),
    .i_Pattern(r_TP_Index),
    .i_HSync(w_HSync_Start),
    .i_VSync(w_VSync_Start),
    .o_HSync(w_HSync_TP),
    .o_VSync(w_VSync_TP),
    .o_Red_Video(w_Red_Video_TP),
    .o_Grn_Video(w_Grn_Video_TP),
    .o_Blu_Video(w_Blu_Video_TP));

    VGA_Sync_Porch #(.VIDEO_WIDTH(c_VIDEO_WIDTH),
                    .TOTAL_COLS(c_TOTAL_COLS),
                    .TOTAL_ROWS(c_TOTAL_ROWS),
                    .ACTIVE_COLS(c_ACTIVE_COLS),
                    .ACTIVE_ROWS(c_ACTIVE_ROWS))
    VGA_Sync_Porch_Inst
    (.i_Clk(i_Clk),
     .i_HSync(w_HSync_TP),
     .i_VSync(w_VSync_TP),
     .i_Red_Video(w_Red_Video_TP),
     .i_Grn_Video(w_Grn_Video_TP),
     .i_Blu_Video(w_Blu_Video_TP),
     .o_HSync(w_HSync_Porch),
     .o_VSync(w_VSync_Porch),
     .o_Red_Video(w_Red_Video_Porch),
     .o_Grn_Video(w_Grn_Video_Porch),
     .o_Blu_Video(w_Blu_Video_Porch));
    
    assign o_VGA_HSync = w_HSync_Porch;
    assign o_VGA_VSync = w_VSync_Porch;

    assign o_VGA_Red_0 = w_Red_Video_Porch[0];
    assign o_VGA_Red_1 = w_Red_Video_Porch[1];
    assign o_VGA_Red_2 = w_Red_Video_Porch[2];
    
    assign o_VGA_Grn_0 = w_Grn_Video_Porch[0];
    assign o_VGA_Grn_1 = w_Grn_Video_Porch[1];
    assign o_VGA_Grn_2 = w_Grn_Video_Porch[2];
    
    assign o_VGA_Blu_0 = w_Blu_Video_Porch[0];
    assign o_VGA_Blu_1 = w_Blu_Video_Porch[1];
    assign o_VGA_Blu_2 = w_Blu_Video_Porch[2];

endmodule